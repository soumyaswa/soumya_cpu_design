`include "mul.sv"
`include "div.sv"
`include "add.sv"
`include "sub.sv"
module top;
  reg [15:0]rs1,rs2;
  wire [15:0]rd,add_rd,co;
  
  reg [3:0]a,b;
  wire [7:0] p;
  
  bit [15:0] greater,equal,less; 
  division dut(rs1,rs2,greater,equal,less); 
  
  //multiplier_4x4 mul_dut(a,b,p);

  //add add_dut(rs1,rs2,add_rd,co);
  //sub sub_dut(rs1,rs2,rd); 
  //mul mul_dut(rs1,rs2,rd);
  //div div_dut(rs1, rs2, rd1,rd2);
 // div div_dut(rs1, rs2, rd);
  initial begin
    repeat(1)begin
      rs1=12;
      rs2=2;
      #1;
      $display("rs1=%d, rs2=%d, greater=%d, equal=%d ,less=%d", rs1,rs2,greater,equal,less); 
     // $display("rs1=%d, rs2=%d, rd=%d", rs1,rs2,rd); 
    //  $display("division output: rs1=%d, rs2=%d, rd1=%d, rd2=%d", rs1,rs2,rd1,rd2); 
      
      /*a=12;
      b=2;
      #5;
      $display("a=%d, b=%d, p=%b", a,b,p);*/
    end
    
  end
  
  initial begin
    $dumpfile("test.vcd");
    $dumpvars(1);
  end
  
endmodule

